LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY sub IS
  GENERIC (
    DATA_WIDTH : INTEGER := 16
  );
  PORT (
    I_1 : IN STD_LOGIC_VECTOR ((DATA_WIDTH - 1) DOWNTO 0);
    I_2 : IN STD_LOGIC_VECTOR ((DATA_WIDTH - 1) DOWNTO 0);
    O : OUT STD_LOGIC_VECTOR ((DATA_WIDTH - 1) DOWNTO 0)
  );
END sub;

ARCHITECTURE Behav OF sub IS
BEGIN
  O <= STD_LOGIC_VECTOR(UNSIGNED(I_2) - UNSIGNED(I_1));
END Behav; -- Behav