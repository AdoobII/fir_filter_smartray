PACKAGE mytypes IS
  TYPE COEFFS IS ARRAY (NATURAL RANGE <>) OF INTEGER;
END PACKAGE;